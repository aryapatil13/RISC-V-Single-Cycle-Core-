`include "pcounter.v"
`include "instruction_memory"

module single_cycle(clk,rst);
   input clk,rst;

endmodule